/home/alexey/tmp/sata2/x393/ddr3/2048Mb_ddr3_parameters.vh