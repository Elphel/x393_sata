/home/alexey/tmp/sata2/x393/ddr3/4096Mb_ddr3_parameters.vh