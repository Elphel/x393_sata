, .INIT_00 (256'h00100000000E0000000C00000033000000200000000A0000000A0000000A0000)
, .INIT_01 (256'h001944521C399446543044170000001900480019040802020204008400220006)
, .INIT_02 (256'h001900050019C82E000C04020090002924FB2502014000190003004204040000)
, .INIT_03 (256'h845284BE44374C682C4214190012003900480018000A01080022001901020050)
, .INIT_04 (256'h00190090003900900019144601020408020202040039B07D707A021000398C6B)
, .INIT_05 (256'h64540C2504580000004E24FB25020420004C24FB25020420005C000000390000)
, .INIT_06 (256'hA47150F8903900600104006B0202003000E2A89368F018E918CB98A758D73882)
, .INIT_07 (256'h0410003900000039B07D00000050004400220039B07D707A307730F000880102)
, .INIT_08 (256'h00050091C88F002200240091288B28FE000C0090008624FB25020140009CD0FB)
, .INIT_09 (256'h48A528A128FE00140039487F0CAD28FE0090009724FB250200C0005004020091)
, .INIT_0A (256'h8839089C020800AD009000AB24FB2502042000500081005048A5002200240039)
, .INIT_0B (256'h00C002080039889C020800090039889C50BA0024002800B5D0FB50F800A000B1)
, .INIT_0C (256'h009000CF24FB250202200039889C50BA00240028009000C5C50224FB24FB0120)
, .INIT_0D (256'h0050C8E028FE000C009000DB24FB25020240003934D2000000D4001100D4C8D2)
, .INIT_0E (256'h00F60082009000ED24FB2502042000390401009000E624FB2502044000500101)
, .INIT_0F (256'h0100020101000021011001000021004400F6000000F6009000F424FB25020420)
, .INIT_10 (256'h0000000000000000000000000000000000000000000000390041000001000000)
, .INITP_00 (256'hC8220098170902401E272722222800309418800820809C802018880022222222)
, .INITP_01 (256'h22082227209C82720A09C22089C680272181A01CB889C8605A2A89C882068270)
, .INITP_02 (256'h0000000000000000000000000000000000000000000000000000000000000082)
