, .INIT_00 (256'h00100000000E0000000C02020035000000220000000C0000000A0000000C0000)
, .INIT_01 (256'h1C3B9448543244190060001B0108001B00500402040401040022000600120000)
, .INIT_02 (256'h001BC8300014000C0210002B24FD25050180001B0003004200180000001B4454)
, .INIT_03 (256'h44394C6A2C44141B0012003B01080028000A04080022001B01020110001B0005)
, .INIT_04 (256'h003B0210001B14480102005004020404003BB07F707C00A0003B8C6D845484C0)
, .INIT_05 (256'h045A0000005024FD25050240004E24FD25050240005E0000003B0000001B0210)
, .INIT_06 (256'h903B02200204006D0402009000E4A89568F218EB18CD98A958D9388464560C27)
, .INIT_07 (256'h0000003BB07F0000005200840022003BB07F707C307930F202080073D10750FA)
, .INIT_08 (256'hC891002200440093288D290100140210008824FD25050180009ED0FF0120003B)
, .INIT_09 (256'h29010024003B48810CAF29010210009924FD250504400052000C009300050093)
, .INIT_0A (256'h003000AF021000AD24FD2505024000520081005248A700220044003B48A728A3)
, .INIT_0B (256'h003B889E00300009003B889E50BC0044008800B7D0FF50FA042000B3883B089E)
, .INIT_0C (256'h24FD25050140003B889E50BC00440048021000C7C50524FD24FD00C000C20030)
, .INIT_0D (256'h29010014021000DD24FD25050280003B34D4000000D6001100D6C8D4021000D1)
, .INIT_0E (256'h021000EF24FD25050240003B0401021000E824FD25050480005201010052C8E2)
, .INIT_0F (256'h002100FF041001030021008400F8000000F8021000F624FD2505024000F80082)
, .INIT_10 (256'h0000000000000000000000000000003B00410107041001030000010302010103)
, .INITP_00 (256'h8220098170902401E272722222800309418810820809C8020188800222222222)
, .INITP_01 (256'h8882227209C82720A09C22089C680272181A01CB889C8605A2A89C882068270C)
, .INITP_02 (256'h0000000000000000000000000000000000000000000000000000000000008888)
