, .INIT_00 (256'h00100000000E0000000C02020035000000220000000C0000000A0000000C0000)
, .INIT_01 (256'h1C3B9448543244190060001B0108001B00500402040401040022000600120000)
, .INIT_02 (256'h001BC8300014000C0210002B2506250D0180001B0003004200180000001B4454)
, .INIT_03 (256'h44394C6A2C44141B0012003B01080028000A04080022001B01020110001B0005)
, .INIT_04 (256'h003B0210001B14480102005004020404003BB07F707C00A0003B8C6D845484C6)
, .INIT_05 (256'h045A000000502506250D0240004E2506250D0240005E0000003B0000001B0210)
, .INIT_06 (256'h903B02200204006D0402009000EDA89868FB18F418D398AF58DF388464560C27)
, .INIT_07 (256'h0000003BB07F0000005200840022003BB07F707C307930FB02080073D10D5103)
, .INIT_08 (256'h0096289029090000000000000014021000882506250D018000A1D1060120003B)
, .INIT_09 (256'h48810CB529090210009C2506250D04400052000C009600050096C89400220044)
, .INIT_0A (256'h024000520081005248AD00220044003B48AD28A929090000000000000024003B)
, .INIT_0B (256'h50C20044008800BDD1065103042000B9883B08A1003000B5021000B32506250D)
, .INIT_0C (256'h00440048021000CDC50D2506250600C000C80030003B88A100300009003B88A1)
, .INIT_0D (256'h0280003B34DA000000DC001100DCC8DA021000D72506250D0140003B88A150C2)
, .INIT_0E (256'h2506250D0480005201010052C8EB29090000000000000014021000E32506250D)
, .INIT_0F (256'h021000FF2506250D024001010082021000F82506250D0240003B0401021000F1)
, .INIT_10 (256'h003B00410410010B0000010B0201010B00210410010B00210084010100000101)
, .INITP_00 (256'h8220098170902401E272722222800309418810820809C8020188800222222222)
, .INITP_01 (256'h89C827209C828009C22089C680272181A01CB889C8605A00AA2722081A00270C)
, .INITP_02 (256'h0000000000000000000000000000000000000000000000000000000020888208)
