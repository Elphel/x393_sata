, .INIT_00 (256'h00100000000E0000000C00000030000000200000000A0000000A0000000A0000)
, .INIT_01 (256'h0019444F1C369443542D44170000001900480019040802020204008400220006)
, .INIT_02 (256'h0019010200500019000C04020090002924F824FF014000190003004204040000)
, .INIT_03 (256'h021000368C68844F84BB44344C652C3F14190012003600480018000A01080022)
, .INIT_04 (256'h00000036000000190090003600900019144301020408020202040036B07A7077)
, .INIT_05 (256'h98A458D4387F64510C2504550000004B24F824FF0420004924F824FF04200059)
, .INIT_06 (256'h30ED008800FFA46E50F590360060010400680202003000DFA89068ED18E618C8)
, .INIT_07 (256'h01400099D0F80410003600000036B07A0000004D004400220036B07A70773074)
, .INIT_08 (256'h004D0402008E0005008EC88C00220024008E288828FB000C0090008324F824FF)
, .INIT_09 (256'h00220024003648A2289E28FB00140036487C0CAA28FB0090009424F824FF00C0)
, .INIT_0A (256'h50F500A000AE88360899020800AA009000A824F824FF0420004D0081004D48A2)
, .INIT_0B (256'h24F824F8012000BD020800368899020800090036889950B70024002800B2D0F8)
, .INIT_0C (256'h001100D1C8CF009000CC24F824FF02200036889950B700240028009000C2C4FF)
, .INIT_0D (256'h0440004D0101004DC8DD28FB000C009000D824F824FF0240003634CF000000D1)
, .INIT_0E (256'h24F824FF042000F30082009000EA24F824FF042000360401009000E324F824FF)
, .INIT_0F (256'h000000FD000000FD020100FD0021011000FD0021004400F3000000F3009000F1)
, .INIT_10 (256'h0000000000000000000000000000000000000000000000000000000000360041)
, .INITP_00 (256'hC3208802605C240900789C9C8888A000C250620020809C802018880022222222)
, .INITP_01 (256'h088820889C827209C828270882271A009C86068072E227218168AA2722081A09)
, .INITP_02 (256'h0000000000000000000000000000000000000000000000000000000000000002)
