, .INIT_00 (256'h00100000000E0000000C00000033000000200000000A0000000A0000000A0000)
, .INIT_01 (256'h001944521C399446543044170000001900880019003002020204008400220006)
, .INIT_02 (256'h001900050019C82E000C04020110002924FB2502024000190003004204040000)
, .INIT_03 (256'h845284BE44374C682C4214190012003900880018000A02080022001901020090)
, .INIT_04 (256'h00190110003901100019144601020030020202040039B07D707A041000398C6B)
, .INIT_05 (256'h64540C2504580000004E24FB250200C0004C24FB250200C0005C000000390000)
, .INIT_06 (256'hA47150F8903900A00104006B0202005000E2A89368F018E918CB98A758D73882)
, .INIT_07 (256'h0060003900000039B07D00000050004400220039B07D707A307730F001080102)
, .INIT_08 (256'h00050091C88F002200240091288B28FE000C0110008624FB25020240009CD0FB)
, .INIT_09 (256'h48A528A128FE00140039487F0CAD28FE0110009724FB25020140005004020091)
, .INIT_0A (256'h8839089C040800AD011000AB24FB250200C000500081005048A5002200240039)
, .INIT_0B (256'h00C004080039889C040800090039889C50BA0024004800B5D0FB50F8012000B1)
, .INIT_0C (256'h011000CF24FB250204200039889C50BA00240028011000C5C50224FB24FB0220)
, .INIT_0D (256'h0050C8E028FE000C011000DB24FB25020440003934D2000000D4001100D4C8D2)
, .INIT_0E (256'h00F60082011000ED24FB250200C000390401011000E624FB2502018000500101)
, .INIT_0F (256'h0100020101000021021001000021004400F6000000F6011000F424FB250200C0)
, .INIT_10 (256'h0000000000000000000000000000000000000000000000390041000001000000)
, .INITP_00 (256'hC8220098170902401E272722222800309418810820809C802018880022222222)
, .INITP_01 (256'h22082227209C82720A09C22089C680272181A01CB889C8605A2A89C882068270)
, .INITP_02 (256'h0000000000000000000000000000000000000000000000000000000000000082)
